///////////////////////////////////
//
//   FILE_NAME   : slave_seq_item.sv
//   Author Name : Ashfaq Manihar
//   Type        : Class
//   Description : 
//   Version     : 1.0
//   Date        : 14/07/2025
//
///////////////////////////////////
`ifndef AXI_SLAVE_SEQ_ITEM_SV
`define AXI_SLAVE_SEQ_ITEM_SV


///////////////////////////////////////////////
/////       WRITE RESPONSE ENUM      //////////
///////////////////////////////////////////////

typedef enum bit[1:0] {
    WRITE_OKAY     = 2'b00,
    WRITE_EXOKAY   = 2'b01,
    WRITE_SLVERR   = 2'b10,
    WRITE_DECERR   = 2'b11 } bresp_en;

///////////////////////////////////////////////
/////       READ RESPONSE ENUM       //////////
///////////////////////////////////////////////

typedef enum bit[1:0] {
    READ_OKAY     = 2'b00,
    READ_EXOKAY   = 2'b01,
    READ_SLVERR   = 2'b10,
    READ_DECERR   = 2'b11 } rresp_en;

///////////////////////////////////////////////
/////       TRANS KIND ENUM          //////////
///////////////////////////////////////////////


typedef enum bit {READ, WRITE} trans_kind_e;

///////////////////////////////////////////////
/////       WRITE BURST ENUM       ////////////
///////////////////////////////////////////////
  
  typedef enum bit[1:0] {
    WRITE_FIXED     = 2'b00,
    WRITE_INCR      = 2'b01,
    WRITE_WRAP      = 2'b10,
    WRITE_RESERVED  = 2'b11 } wburst_en;

///////////////////////////////////////////////
/////       READ BURST ENUM        ////////////
///////////////////////////////////////////////

  typedef enum bit[1:0] {
    READ_FIXED     = 2'b00,
    READ_INCR      = 2'b01,
    READ_WRAP      = 2'b10,
    READ_RESERVED  = 2'b11 } rburst_en;

///////////////////////////////////////////////
/////       WRITE SIZE ENUM        ////////////
///////////////////////////////////////////////

typedef enum bit[2:0] {
    WRITE_1_BYTE     = 3'b000,
    WRITE_2_BYTE     = 3'b001,
    WRITE_4_BYTE     = 3'b010,
    WRITE_8_BYTE     = 3'b011,  
    WRITE_16_BYTE      = 3'b100,
    WRITE_32_BYTE      = 3'b101,
    WRITE_64_BYTE      = 3'b110,
    WRITE_128_BYTE     = 3'b111 } wsize_en;


///////////////////////////////////////////////
/////       READ SIZE ENUM         ////////////
///////////////////////////////////////////////

typedef enum bit[2:0] {
    READ_1_BYTE     = 3'b000,
    READ_2_BYTE     = 3'b001,
    READ_4_BYTE     = 3'b010,
    READ_8_BYTE     = 3'b011,  
    READ_16_BYTE    = 3'b100,
    READ_32_BYTE    = 3'b101,
    READ_64_BYTE    = 3'b110,
    READ_128_BYTE   = 3'b111 } rsize_en;



class slave_seq_item #(parameter ADDR_WIDTH = 32,DATA_WIDTH =32) extends uvm_sequence_item;
  
  trans_kind_e kind;
   
  // Write Address Channel
   bit [7:0]              AWID;
   bit [ADDR_WIDTH-1:0]   AWADDR[$];   // QUEUE to store further transfers address 
   bit [7:0]              AWLEN;
   wsize_en               AWSIZE;
   wburst_en              AWBURST;


  // Write Data Channel
   bit [7:0]              WID;
   bit [DATA_WIDTH-1:0]   WDATA[$];       //To store data from the master driver
   rand bit [DATA_WIDTH/8-1:0] WSTRB[$];    //THINK: whether the WSTRB should be generated by the slave or the interconect ?


  // Write Response Channel
  rand bit [7:0]          BID;
  bresp_en                BRESP;


  // Read Address Channel
  bit [7:0]              ARID;
  bit [ADDR_WIDTH-1:0]   ARADDR[$];       // QUEUE to store further read address 

  bit [7:0]              ARLEN;
  rsize_en               ARSIZE;
  rburst_en              ARBURST;


  // Read Data Channel
  rand bit [7:0]              RID;
  rand bit [DATA_WIDTH-1:0]   RDATA[$];
  rresp_en                    RRESP;


       
  `uvm_object_param_utils_begin(slave_seq_item #(ADDR_WIDTH, DATA_WIDTH))
//     `uvm_field_enum(trans_type_e, trans_type, UVM_ALL_ON)

    `uvm_field_int(AWID,      UVM_ALL_ON)
    `uvm_field_queue_int(AWADDR, UVM_ALL_ON)
    `uvm_field_int(AWLEN,     UVM_ALL_ON)
    `uvm_field_enum(wburst_en, AWBURST , UVM_ALL_ON)
    `uvm_field_enum(trans_kind_e, kind, UVM_ALL_ON)
    `uvm_field_int(WID,      UVM_ALL_ON)

    `uvm_field_queue_int(WDATA, UVM_ALL_ON)
    `uvm_field_queue_int(WSTRB,     UVM_ALL_ON)    
    `uvm_field_enum(wsize_en, AWSIZE, UVM_ALL_ON)

    `uvm_field_int(ARID,      UVM_ALL_ON)
   `uvm_field_queue_int(ARADDR, UVM_ALL_ON)
    `uvm_field_enum(rsize_en, ARSIZE, UVM_ALL_ON)   
    `uvm_field_int(ARLEN,     UVM_ALL_ON)
    `uvm_field_enum(rburst_en, ARBURST , UVM_ALL_ON)
    `uvm_field_queue_int(RDATA, UVM_ALL_ON) 
    `uvm_field_int(RID,       UVM_ALL_ON)

  `uvm_object_utils_end



 
  
  function new(string name = "slave_seq_item");
    super.new(name);
  endfunction
  
endclass

`endif


